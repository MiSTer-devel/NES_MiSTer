module MicroCodeTableInner
(
	input clk,
	input ce,
	input reset,
	input [7:0] IR,
	input [2:0] State,
	output reg [8:0] M
);

wire [8:0] L[2048] = '{
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_10_10100, // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
	9'b00_10_10100, // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
	9'b00_10_10101, // P->[SP--]
	9'b00_11_00011, // [VECT]->T
	9'b10_11_10011, // [VECT]:T->PC
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00011, // [PC]->
	9'b10_10_01111, // P->[SP--]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_10_10100, // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
	9'b00_10_10100, // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
	9'b00_10_00111, // KEEP_AC
	9'b10_00_10011, // [PC]:T->PC
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00011, // [PC]->
	9'b00_10_10000, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	9'b10_10_00010, // ['ALU([SP])->A', '[SP]->P']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_10_10000, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	9'b00_10_10110, // [SP]->P,SP+1->SP
	9'b00_10_10000, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	9'b10_10_10011, // [SP]:T->PC
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00011, // [PC]->
	9'b10_10_01110, // ALU(A)->[SP--]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_00_10011, // [PC]:T->PC
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_10_10000, // SP+1->SP
	9'bxx_xx_xxxxx, // []
	9'b00_10_10000, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	9'b00_10_10011, // [SP]:T->PC
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00011, // [PC]->
	9'b00_10_10000, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	9'b10_10_00010, // ['ALU([SP])->A', '[SP]->P']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00001, // [PC++]->AH
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b10_01_10011, // [AX]:T->PC
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_10010, // X->S
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00110, // ALU()->[AX]
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_00111, // [AX]->?,AL+X->AL
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01011, // [AX]->AH,T->AL
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00000, // ['[PC++]->AL', '[PC++]->T']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_01101, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_00001, // [PC++]->AH
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00000, // ['[PC++]->?', 'PC+1->PC', '']
	9'b11_00_10001, // PC+T->PC
	9'bxx_xx_xxxxx, // []
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b01_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_01_01010, // [AX]->T,AL+1->AL
	9'b00_01_01100, // [AX]->AH,T+Y->AL
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_01_00111, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00010, // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->X,Y', 'ALU()->A']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b10_00_00011, // ['NO-OP', '']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00011, // ['ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b01_00_01000, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b10_01_00010, // ['ALU([AX])->A', 'ALU([AX])->?']
	9'bxx_xx_xxxxx, // []
	9'bxx_xx_xxxxx, // []
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101, // T->[AX]
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b00_00_00000, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
	9'b11_00_01000, // ['[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+Y->AL']
	9'bxx_xx_xxxxx, // []
	9'b00_01_01001, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	9'b00_01_00011, // [AX]->T
	9'b00_01_00100, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	9'b10_01_00101  // T->[AX]
};

always @(posedge clk) begin
	if (reset) begin
		M <= 0; // Stupid XILINX inferral only allows 0 as reset value.
	end else if (ce) begin
		M <= L[{IR, State}];    
	end
end

endmodule

module MicroCodeTable
(
	input clk,
	input ce,
	input reset,
	input [7:0] IR,
	input [2:0] State,
	output [37:0] Mout
);

wire [8:0] M;
MicroCodeTableInner inner
(
	clk,
	ce,
	reset,
	IR,
	State, M
);

wire [14:0] A[32] = '{
	15'b_10__0_10101_0xx_01_00, // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T', 'PC+1->PC', '']
	15'b_xx__0_0xx11_0xx_01_00, // [PC++]->AH
	15'b_xx__1_00000_0xx_00_00, // ['ALU([AX])->A', 'ALU([AX])->?', '[PC]->,ALU()->A', 'Setappropriateflags', 'ALU([SP])->A', '[SP]->P', 'ALU()->X,Y', 'ALU()->A']
	15'b_10__0_00000_0xx_00_00, // ['[AX]->T', 'ALU([AX])->?', 'ALU([AX])->A', 'ALU([AX])->', '[PC]->', 'NO-OP', '[VECT]->T', '']
	15'b_11__1_00000_100_00_00, // ['T->[AX],ALU(T)->T', 'T->[AX],ALU(T)->T:A']
	15'b_xx__0_xxxxx_100_00_00, // T->[AX]
	15'b_xx__0_00000_101_00_00, // ALU()->[AX]
	15'b_0x__0_10000_0xx_00_00, // ['[AX]->?,AL+X->AL', '[AX]->?,AL+X/Y->AL', 'KEEP_AC']
	15'b_xx__0_10011_0xx_01_00, // ['[PC++]->AH,AL+X/Y->AL', '[PC++]->AH,AL+X->AL', '[PC++]->AH,AL+Y->AL']
	15'b_10__0_0xx10_0xx_00_00, // ['[AX]->?,AH+FIX->AH', '[AX]->T,AH+FIX->AH']
	15'b_10__0_11000_0xx_00_00, // [AX]->T,AL+1->AL
	15'b_xx__0_11111_0xx_00_00, // [AX]->AH,T->AL
	15'b_xx__0_10011_0xx_00_00, // [AX]->AH,T+Y->AL
	15'b_xx__1_xxxxx_0xx_01_00, // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
	15'b_xx__0_xxxxx_101_00_11, // ALU(A)->[SP--]
	15'b_xx__0_xxxxx_110_00_11, // P->[SP--]
	15'b_10__0_xxxxx_0xx_00_10, // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
	15'b_xx__0_xxxxx_0xx_11_00, // PC+T->PC
	15'b_xx__0_xxxxx_0xx_00_01, // X->S
	15'b_xx__0_xxxxx_0xx_10_00, // ['[PC]:T->PC', '[AX]:T->PC', '[VECT]:T->PC', '[SP]:T->PC']
	15'b_0x__0_xxxxx_111_00_11, // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
	15'b_xx__1_xxxxx_110_00_11, // P->[SP--]
	15'b_xx__1_xxxxx_0xx_00_10, // [SP]->P,SP+1->SP
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx, // []
	15'b_xx__x_xxxxx_xxx_xx_xx  // []
};

wire [18:0] B[256] = '{
	19'bxxxxxxxxxx0_000_00_010, 19'b000010x0001_010_00_001, 19'bxx0100010x0_000_00_001, 19'b00010000001_010_00_001, 
	19'b000010x0000_xxx_00_xxx, 19'b000010x0001_010_00_001, 19'bxx0100010x0_000_00_001, 19'b00010000001_010_00_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0001_010_00_001, 19'b001000010x0_010_00_001, 19'b000010x0001_010_00_001, 
	19'b000010x0000_xxx_00_xxx, 19'b000010x0001_010_00_001, 19'bxx0100010x0_000_00_001, 19'b00010000001_010_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x0001_010_11_001, 19'bxx0100010x0_000_11_001, 19'b00010000001_010_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0001_010_00_001, 19'bxx0100010x0_000_00_001, 19'b00010000001_010_00_001, 
	19'bxxxxxxxxxx0_000_10_101, 19'b000010x0001_010_10_001, 19'bxx0100010x0_000_10_001, 19'b00010000001_010_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0001_010_00_001, 19'bxx0100010x0_000_00_001, 19'b00010000001_010_00_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0011_010_00_001, 19'bxx0100110x0_000_00_001, 19'b00010010011_010_00_001, 
	19'b000010x0010_000_00_001, 19'b000010x0011_010_00_001, 19'bxx0100110x0_000_00_001, 19'b00010010011_010_00_001, 
	19'bxxxxxxxxxx0_000_00_100, 19'b000010x0011_010_00_001, 19'b001000110x0_010_00_001, 19'b000010x0011_010_00_001, 
	19'b000010x0010_000_00_001, 19'b000010x0011_010_00_001, 19'bxx0100110x0_000_00_001, 19'b00010010011_010_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x0011_010_11_001, 19'bxx0100110x0_000_11_001, 19'b00010010011_010_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0011_010_00_001, 19'bxx0100110x0_000_00_001, 19'b00010010011_010_00_001, 
	19'bxxxxxxxxxx0_000_10_101, 19'b000010x0011_010_10_001, 19'bxx0100110x0_000_10_001, 19'b00010010011_010_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0011_010_00_001, 19'bxx0100110x0_000_00_001, 19'b00010010011_010_00_001, 
	19'bxxxxxxxxxx0_000_00_100, 19'b000010x0101_010_00_001, 19'bxx0101010x0_000_00_001, 19'b00010100101_010_00_001, 
	19'b000010x0100_xxx_00_xxx, 19'b000010x0101_010_00_001, 19'bxx0101010x0_000_00_001, 19'b00010100101_010_00_001, 
	19'b001010x10x0_xxx_00_xxx, 19'b000010x0101_010_00_001, 19'b001001010x0_010_00_001, 19'b000010x0101_010_00_001, 
	19'bxxxxxxxxxx0_000_00_001, 19'b000010x0101_010_00_001, 19'bxx0101010x0_000_00_001, 19'b00010100101_010_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x0101_010_11_001, 19'bxx0101010x0_000_11_001, 19'b00010100101_010_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0101_010_00_001, 19'bxx0101010x0_000_00_001, 19'b00010100101_010_00_001, 
	19'bxxxxxxxxxx0_000_10_110, 19'b000010x0101_010_10_001, 19'bxx0101010x0_000_10_001, 19'b00010100101_010_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0101_010_00_001, 19'bxx0101010x0_000_00_001, 19'b00010100101_010_00_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0111_010_00_001, 19'bxx0101110x0_000_00_001, 19'b00010110111_010_00_001, 
	19'b000010x0110_xxx_00_xxx, 19'b000010x0111_010_00_001, 19'bxx0101110x0_000_00_001, 19'b00010110111_010_00_001, 
	19'bxx0010x10x0_010_00_001, 19'b000010x0111_010_00_001, 19'b001001110x0_010_00_001, 19'b000010x0111_010_00_001, 
	19'bxxxxxxxxxx0_000_00_001, 19'b000010x0111_010_00_001, 19'bxx0101110x0_000_00_001, 19'b00010110111_010_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x0111_010_11_001, 19'bxx0101110x0_000_11_001, 19'b00010110111_010_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0111_010_00_001, 19'bxx0101110x0_000_00_001, 19'b00010110111_010_00_001, 
	19'bxxxxxxxxxx0_000_10_110, 19'b000010x0111_010_10_001, 19'bxx0101110x0_000_10_001, 19'b00010110111_010_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x0111_010_00_001, 19'bxx0101110x0_000_00_001, 19'b00010110111_010_00_001, 
	19'b011010x10x0_xxx_00_xxx, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_xxx_00_xxx, 19'b111010x10x1_xxx_00_xxx, 
	19'b011010x10x0_xxx_00_xxx, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_xxx_00_xxx, 19'b111010x10x1_xxx_00_xxx, 
	19'b011011010x0_100_00_001, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_010_00_001, 19'b111010x10x1_xxx_00_xxx, 
	19'b011010x10x0_xxx_00_xxx, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_xxx_00_xxx, 19'b111010x10x1_xxx_00_xxx, 
	19'b011010x10x0_xxx_11_xxx, 19'b001010x10x1_xxx_11_xxx, 19'b101010x10x0_xxx_11_xxx, 19'b111010x10x1_xxx_11_xxx, 
	19'b011010x10x0_xxx_00_xxx, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_xxx_10_xxx, 19'b111010x10x1_xxx_10_xxx, 
	19'b011010x10x0_010_10_001, 19'b001010x10x1_xxx_10_xxx, 19'b101010x10x0_xxx_10_xxx, 19'b111010x10x1_xxx_10_xxx, 
	19'b011010x10x0_xxx_00_xxx, 19'b001010x10x1_xxx_00_xxx, 19'b101010x10x0_xxx_10_xxx, 19'b111010x10x1_xxx_10_xxx, 
	19'bxx0010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'bxx0010x10x0_001_00_001, 19'bxx0010x10x1_011_00_001, 
	19'bxx0010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'bxx0010x10x0_001_00_001, 19'bxx0010x10x1_011_00_001, 
	19'b001010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'b001010x10x0_001_00_001, 19'bxx0010x10x1_011_00_001, 
	19'bxx0010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'bxx0010x10x0_001_00_001, 19'bxx0010x10x1_011_00_001, 
	19'bxx0010x10x0_xxx_11_xxx, 19'bxx0010x10x1_010_11_001, 19'bxx0010x10x0_xxx_11_xxx, 19'bxx0010x10x1_011_11_001, 
	19'bxx0010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'bxx0010x10x0_001_10_001, 19'bxx0010x10x1_011_10_001, 
	19'bxx1110x10x0_000_10_011, 19'bxx0010x10x1_010_10_001, 19'bxx1110x10x0_001_10_001, 19'bxx0010x10x1_xxx_10_xxx, 
	19'bxx0010x10x0_100_00_001, 19'bxx0010x10x1_010_00_001, 19'bxx0010x10x0_001_10_001, 19'bxx0010x10x1_011_10_001, 
	19'b010010x1100_000_00_001, 19'b000010x1101_000_00_001, 19'bxx0111010x0_000_00_001, 19'b00011101101_000_00_001, 
	19'b010010x1100_000_00_001, 19'b000010x1101_000_00_001, 19'bxx0111010x0_000_00_001, 19'b00011101101_000_00_001, 
	19'b011011110x0_100_00_001, 19'b000010x1101_000_00_001, 19'b101011010x0_001_00_001, 19'b000010x1101_000_00_001, 
	19'b010010x1100_000_00_001, 19'b000010x1101_000_00_001, 19'bxx0111010x0_000_00_001, 19'b00011101101_000_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x1101_000_11_001, 19'bxx0111010x0_000_11_001, 19'b00011101101_000_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x1101_000_00_001, 19'bxx0111010x0_000_00_001, 19'b00011101101_000_00_001, 
	19'bxxxxxxxxxx0_000_10_111, 19'b000010x1101_000_10_001, 19'bxx0111010x0_000_10_001, 19'b00011101101_000_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x1101_000_00_001, 19'bxx0111010x0_000_00_001, 19'b00011101101_000_00_001, 
	19'b100010x1100_000_00_001, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b00011111111_010_00_001, 
	19'b100010x1100_000_00_001, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b00011111111_010_00_001, 
	19'b101011110x0_001_00_001, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b000010x1111_010_00_001, 
	19'b100010x1100_000_00_001, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b00011111111_010_00_001, 
	19'bxxxxxxxxxx0_xxx_11_xxx, 19'b000010x1111_010_11_001, 19'bxx0111110x0_000_11_001, 19'b00011111111_010_11_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b00011111111_010_00_001, 
	19'bxxxxxxxxxx0_000_10_111, 19'b000010x1111_010_10_001, 19'bxx0111110x0_000_10_001, 19'b00011111111_010_10_001, 
	19'bxxxxxxxxxx0_xxx_00_xxx, 19'b000010x1111_010_00_001, 19'bxx0111110x0_000_00_001, 19'b00011111111_010_00_001
};

wire [14:0] R = A[M[4:0]];
reg [18:0] AluFlags;
always @(posedge clk) begin
	if (reset) begin
		AluFlags <= 0;
	end else if (ce) begin  
		AluFlags <= B[IR];
	end
end

assign Mout = {
	AluFlags,// 19
	M[8:7],  // NextState // 2
	R[14:13],// LoadT     // 2
	R[12],   // FlagCtrl  // 1
	R[11:7], // AddrCtrl  // 5
	R[6:4],  // MemWrite  // 3
	M[6:5],  // AddrBus   // 2
	R[3:2],  // LoadPC    // 2
	R[1:0]   // LoadSP    // 2
};

endmodule

